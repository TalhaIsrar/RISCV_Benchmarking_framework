module if_id_pipeline(
    input clk,
    input rst,
    input pipeline_flush,
    input pipeline_en,
        
    input if_flush,
    input [31:0] if_pc,
    input [31:0] if_instruction,
    input if_pred_taken,
    input if_pred_valid,
    input [31:0] if_predicted_pc,

    output reg id_flush,
    output reg [31:0] id_pc,
    output [31:0] id_instruction,
    output reg [31:0] id_predicted_pc,
    output reg id_pred_taken,
    output reg id_pred_valid
);

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            id_pc <= 32'h00000000;
            id_pred_taken <= 1'b0;
            id_flush <= 1'b0;
            id_predicted_pc <= 0;
            id_pred_valid <= 0;
        end else if (pipeline_flush) begin
            id_pc <= id_pc;
            id_pred_taken <= 1'b0;
            id_flush <= if_flush;
            id_predicted_pc <= 0;
            id_pred_valid <= 0;
        end else if (pipeline_en) begin
            id_pc <= if_pc;
            id_pred_taken <= if_pred_taken;  
            id_flush <= if_flush; 
            id_predicted_pc <= if_predicted_pc;
            id_pred_valid <= if_pred_valid;
        end
    end

    // Instruction is passed directly from fetch stage to decode stage because
    // register already in instruction memory module
    assign id_instruction = if_instruction;

endmodule