module fetch_stage(
    input logic clk,
    input logic rst,
    input logic pc_en,
    input logic flush,
    input logic [31:0] pc_jump_addr,
    input logic jump_en,
    input logic [31:0] btb_target_pc,
    input logic btb_pc_valid,
    input logic btb_pc_predictTaken,
    output logic [31:0] instruction,
    output logic [31:0] pc
);
    
    wire [31:0] next_pc;

    // Instantiate the PC module
    pc pc_inst (
        .clk(clk),
        .rst(rst),
        .next_pc(next_pc),
        .pc_en(pc_en),
        .pc(pc)
    );

    // Instantiate the PC update module
    pc_update pc_update_inst (
        .pc(pc),
        .pc_jump_addr(pc_jump_addr),
        .btb_target_pc(btb_target_pc),
        .btb_pc_valid(btb_pc_valid),
        .btb_pc_predictTaken(btb_pc_predictTaken),
        .jump_en(jump_en),
        .next_pc(next_pc)
    );

    // Instantiate the instruction memory module
    instruction_mem instruction_mem_inst (
        .clk(clk),
        .rst(rst),
        .pc(pc),
        .read_en(pc_en),
        .write_en(1'b0),
        .flush(flush),
        .write_addr(14'd0),
        .write_data(32'h00000000),
        .instruction(instruction)
    );

endmodule